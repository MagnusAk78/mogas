signIn = Logga in
signUp = Registrera dig
signOut = Logga ut

language = Språk
welcome = Välkommen {0}
welcomeLeadMessage = Det här är en webb applikation som kan hjälpa er att administrera ett automationssystem.
welcomeInfoMessage = Börja med att skapa en domän (organisation/system/fabrik). Navigera dig fram i navigationsrutan till höger eller högst upp under bläddra.
diveIn = Börja

firstName = Förnamn
lastName = Efternman
name = Namn
email = Epost
password = Lösenord
rememberMe = Kom ihåg mig
shortText = Kort text
text = Text

activeDomain = Aktiv domän: {0}
noActiveDomain = Ingen aktiv domän

navigation = Navigera
list = Lista
create = Skapa ny
domains = Domäner
users = Användare
browse = Bläddra
instructions = Instruktioner
issues = Avvikelser

createDomain = Skapa ny domän
amlFiles = AML filer
parseAmlFiles = Generera databas
uploadAmlFile = Ladda upp AML fil
image = Bild
video = Video
changeImage = Byt bild
manageUsers = Hantera användare
chooseActiveDomain = Välj aktiv domän
rearrange = Omarrangera

details = Detaljer
newInstruction = Ny instruktion
newIssue = Ny avvikelse
addMore = Lägg till fler
addTo = Addera till {0}

editAllowedUsers = Tillåtna användare för {0}
thereMustBeAtLeastOneAllowedUser = Det måste finnas minst en användare

edit = Editera: {0}
delete = Ta bort

fileRemoved = Fil bortplockad

chooseImageFile = Välj bild fil
imageUpload = Ladda upp bild