command.new = Ny
command.add = Lägg till
command.update = Uppdatera
command.delete = Ta bort
command.edit = Editera
command.back = Tillbaka
command.previous = Föregående
command.next = Nästa
command.go.back = Gå tillbaka
command.go.further = Gå vidare

navigation.organisations = Org.
navigation.users = Anv.
navigation.factories = Bläddra
navigation.instructions = Instr.
navigation.issues = Avvikelser

home = Välkommen
home.welcome = Välkommen {0} {1}

language = Språk

link.video = Se film

function.list = Lista
function.create = Skapa ny
function.edit = Ändra
function.details = Detaljer

organisations = Organisationer
organisation.name = Organisationsnamn
organisation.allowedUsers = Godkända användare
organisation.changeAllowedUsers = Editera godkända användare
organisation.minimum.one.user = Det måste finnas minst en godkänd användare
organisations.select.active = Välj aktiv organisation
organisations.active.organisation = Aktiv organisation
organisation.remove.self.not.allowed = Det är inte tillåtet att ta bort inloggad användare

users = Användare
user.details = Info om användare
user.username = Användarnamn
user.password = Lösenord
user.confirmPassword = Bekräfta lösenord
user.firstName = Förnamn
user.lastName = Efternamn
user.email = epost
user.active.organisation = Aktiv organisation
user.editAccount = Editera användaruppgifter
user.signOut = Logga ut
user.signIn = Logga in
user.signUp = Registrera konto
user.question.notMember = Ej registrerad?
user.question.alreadyMember = Redan registrerad?
user.allowed.organisations = Tillåtna organisationer

factories = Fabriker
factory.view.hierarchy = Se fabriksträd
factory.hierarchy = Fabriksträd {0}
factory.hierarchies = Fabriksträd
factory.element = Fabrikselement: {0}
factory.element.ie = Fabrikselement
factory.element.ei = Extern koppling/interface
factory.add.amlfile = Lägg till AML-fil
factory.add.image = Lägg till bildfil

instructions = Instruktioner
instruction = Instruktion
instruction.create = Skapa instruktion
instruction.title = Titel
instruction.textDescription = Beskrivning
instruction.refers.to = Avser: {0}
instruction.show.created.by = Skapad av {0}
instruction.orderNumber = nummer
instruction.show.orderNumber = nr: {0}
instruction.show.created.by = Skapad av {0}
instructions.show = Instruktioner

instructions.move.down = Flytta ner
instructions.move.up = Flytta upp

issues = Avvikelser
issue = Avvikelse
issue.create = Skapa avvikelse
issue.title = Titel
issue.textDescription = Beskrivning
issue.assignedTo = Tilldelad användare
issue.priority = Prioritet
issues.list.all = Alla avvikelser
issues.list.all.open = Öppna avvikelser
issues.list.all.my.open = Mina öppna avvikelser
issue.close = Stäng denna avvikelse
issue.reopen = Återöppna
issue.refers.to = Avser: {0}

issue.show.priority = Prioritet: {0}
issue.show.not.assigned = Inte tilldelad någon användare
issue.show.assigned.to = Tilldelad {0}
issue.show.open = Öppen
issue.show.closed = Stängd
issue.show.created.by = Skapad av {0}
issue.show.history = Historik

issue.create.new = Rapportera avvikelse

AmlHierarchy.name = {0} (Hierarkinamn)
ExternalInterface = EI {0}
InternalElement = IE {0}

image.file = Bild

validation.duplicate = Dubblett

db.success.save = {0} skapad
db.success.remove = {0} borttagen
db.success.update = {0} uppdaterad

db.error.write = Problem att spara till databas
db.error.read = Problem att läsa från databas
db.error.find = Hittade inte {0}:{1} i databas
db.error.dependencies = Det finns beroenden (minst till {0})
db.error.read.file = Fel vid läsning av fil: {0}
db.error.missing = {0} verkar inte finnas

upload.error.notAllowedContentType = Filen är inte av tillåten typ (mime/content-type)

signupVerification.passwords.doNotMatch = Lösenorden matchar inte
signupVerification.email.taken = Det finns redan en användare med detta epostaddress
signupVerification.username.taken = Det finns redan en användare med detta användarnamn

invalid.credentials = Fel användarnamn eller lösenord
access.denied = Icke behörig
not.set = Inte valt
select.active.organisation = Välj aktiv organisation
upload.image = Ladda upp bild
change.upload.image = Byt/ladda up bild
no.assigned.user = [Inte tilldedad]
none = ingen